library IEEE;
use IEEE.std_logic_1164.all;

entity sumresNb_tb is
end;

architecture sumresNb_tb_arq of sumresNb_tb is
	
	constant N_tb: natural := 4;
	
	-- Declaracion de senales de prueba
	signal a_tb: std_logic_vector(N_tb-1 downto 0) := (N_tb-1 downto 0 => '0');
	signal b_tb: std_logic_vector(N_tb-1 downto 0) := (N_tb-1 downto 0 => '0');
	signal ci_tb: std_logic := '0';
	signal s_tb: std_logic_vector(N_tb-1 downto 0);
	signal co_tb: std_logic;

begin

	a_tb <=  "0111" after 100 ns, "1000" after 300 ns,"1100" after 500 ns;
	b_tb <=  "0100" after 200 ns, "0011" after 400 ns,"0010" after 600 ns;
	ci_tb <= not ci_tb after 50 ns;

	DUT: entity work.sumresNb
		generic map(
			N => N_tb
		)
		port map(
			a_i	 => a_tb, 
			b_i	 => b_tb,
			ci_i => ci_tb,
			s_o	 => s_tb,
			co_o => co_tb
		);
	
end;